      	
parameter first = 8'b0000_0001, second = 8'b0000_0010,third = 8'b0000_0100, fourth = 8'b0000_1000, fifth = 8'b0001_0000,sixth=8'b0010_0000,seventh=8'b0100_0000,eighth=8'b1000_0000;	
